`ifndef COMP_DONE
`define COMP_DONE

package definitions;

	parameter VERSION="1.0a";
	parameter ENGINEER="Diego HR";

endpackage

import definitions::*;

`endif